library verilog;
use verilog.vl_types.all;
entity top is
    port(
        inputs          : in     vl_logic;
        real_out        : out    vl_logic
    );
end top;
